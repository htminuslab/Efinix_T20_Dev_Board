---------------------------------------------------------------------------------------------------
--                                                                           
--  T20Q100 Simple PLL test, toggle LED with a 48MHz clock
--                                         
--  Copyright (C) 2025 HT-LAB                                           
--                                                                                                            
--  https://github.com/htminuslab    
--                                                                             
---------------------------------------------------------------------------------------------------        
--
--  Simple test to toggle the 3 LED's, the clock is 48MHz generated by a PLL
--  
--
--
--  Revision History:                                                        
--                                                                           
--  Date:          Revision         Author         
--  14-jun-2025	   1.0				HABT
---------------------------------------------------------------------------------------------------
library IEEE;
use IEEE.std_logic_1164.all;
use ieee.numeric_std.all;

entity plltest is
	port (	RESETN	: in  std_logic;
			CLK		: in  std_logic;
			LED1   	: out std_logic;
			LED2   	: out std_logic;
			LED3   	: out std_logic);
end plltest;

architecture rtl of plltest is

	component EFX_PLL_V2 is
	generic ( N, M, O        : integer := 1;
			  CLKOUT0_DIV    : integer := 1;
			  CLKOUT1_DIV    : integer := 1;
			  CLKOUT2_DIV    : integer := 1;
			  CLKOUT0_PHASE  : integer := 0;
			  CLKOUT1_PHASE  : integer := 0;
			  CLKOUT2_PHASE  : integer := 0;
			  FEEDBACK_CLK   : string := "INTERNAL";
			  FEEDBACK_MODE  : string := "INTERNAL";
			  REFCLK_FREQ    : real := 25.0);
	port ( CLKOUT0, CLKOUT1, CLKOUT2, LOCKED : out std_logic;
		   RSTN, FBK                         : in  std_logic;
		   CLKIN                             : in  std_logic_vector(3 downto 0);
		   CLKSEL                            : in  std_logic_vector(1 downto 0));
	end component EFX_PLL_V2;

	signal CLKOUT0_s   : std_logic;
	signal counter  : unsigned(25 downto 0);		-- divide 48MHz

begin

    ----------------------------------------------------
    -- PLL Instantiation, requires Unified netlist mode
    ----------------------------------------------------
	EFX_PLL_V2_inst : EFX_PLL_V2					
	generic map (
		M => 128,
		N => 1,
		O => 2,
		CLKOUT0_DIV   => 8,
		CLKOUT1_DIV   => 2,
		CLKOUT2_DIV   => 2,
		CLKOUT0_PHASE => 0,
		CLKOUT1_PHASE => 0,
		CLKOUT2_PHASE => 0,
		FEEDBACK_CLK  => "INTERNAL",
		FEEDBACK_MODE => "INTERNAL",
		REFCLK_FREQ   => 12.0
	)
	port map (
		CLKOUT0 => CLKOUT0_s,             
		CLKOUT1 => open,
		CLKOUT2 => open,
		LOCKED  => open,
		RSTN    => RESETN,
		FBK     => '0',
		CLKIN   => "000"&CLK,
		CLKSEL  => "00"
	);

    process (CLKOUT0_s,RESETN)
	begin
		if RESETN='0' then
			counter  <= (others => '0');
		elsif rising_edge(CLKOUT0_s) then
			counter <= counter+1;
		end if;
	end process;
	    
    LED1 <= counter(23);	
	LED2 <= counter(24);
	LED3 <= counter(25);

end rtl;
