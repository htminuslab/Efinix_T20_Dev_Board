---------------------------------------------------------------------------------------------------
--                                                                           
--  T20Q100 Led toggle test
--                                         
--  Copyright (C) 2025 HT-LAB                                           
--                                                                                                            
--  https://github.com/htminuslab    
--                                                                             
---------------------------------------------------------------------------------------------------        
--
--  Simple test to toggle the 3 LED's, the clock is 12MHz generated by the STMC071
--  
--
--
--  Revision History:                                                        
--                                                                           
--  Date:          Revision         Author         
--  14-jun-2025	   1.0				HABT
---------------------------------------------------------------------------------------------------
library IEEE;
use IEEE.std_logic_1164.all;
use ieee.numeric_std.all;

entity blink is
	port (	RESETN	: in  std_logic;
			CLK		: in  std_logic;
			LED1   	: out std_logic;
			LED2   	: out std_logic;
			LED3   	: out std_logic);
end blink;

architecture rtl of blink is

	signal counter  : unsigned(23 downto 0);		-- 12MHz, 1 sec=B71B00 5B8D80

begin

    process (CLK,RESETN)
	begin
		if RESETN='0' then
			counter  <= (others => '0');
		elsif rising_edge(CLK) then
			counter <= counter+1;
		end if;
	end process;
	    
    LED1 <= counter(21);	
	LED2 <= counter(22);
	LED3 <= counter(23);

end rtl;
